**********************************
* xor_fakeNMOS test netlist
**********************************
.option post=2 
.lib sm046005-1j.hspice typical
.param Wp=2um Wn=1um dd=3.3V cf=0.1PF NL=0.35um PL=0.35um
.global VDD GND

.subckt cmos_inv IN Y_inv
MN   Y_inv   IN    GND   GND   NMOS_3P3   W=Wn  L=0.35um
MP   Y_inv   IN    VDD   VDD   PMOS_3P3   W=Wp  L=0.35um
.ENDS

* NMOS: D G S SUB 
* PMOS: D G S SUB

* .subckt AND2 A B Y_inv
* N1   a       B    GND   GND   NMOS_3P3   W=Wn   L=NL
* N2   Y_inv   A    a     a     NMOS_3P3   W=Wn   L=NL
* P1   Y_inv   A    VDD   VDD   PMOS_3P3   W=Wp   L=PL
* P2   Y_inv   B    VDD   VDD   PMOS_3P3   W=Wp   L=PL   
* .ends

.subckt AND2 IN1 IN2 Y
MN1   a       IN2    GND   GND   NMOS_3P3   W=2*Wn   L=0.35um
MN2   Y_inv   IN1    a     a     NMOS_3P3   W=2*Wn   L=0.35um
MP1   Y_inv   IN1    VDD   VDD   PMOS_3P3   W=Wp   L=0.35um
MP2   Y_inv   IN2    VDD   VDD   PMOS_3P3   W=Wp   L=0.35um 

MN3   Y       Y_inv  GND   GND   NMOS_3P3   W=Wn   L=0.35um
MP3   Y       Y_inv  VDD   VDD   PMOS_3P3   W=Wp   L=0.35um
.ends


X1 A0 B0 Y AND2
* X2 Y_inv Y cmos_inv

* X1 A A1 VDD GND cmos_inv
* X2 B B1 VDD GND cmos_inv
* MN1   A1  B1    Y   GND   NMOS_3P3   W=1um L=0.35um
* MP1   A1  B     Y   VDD   PMOS_3P3   W=Wp  L=0.35um
* MN2   A   B     Y   GND   NMOS_3P3   W=1um L=0.35um
* MP2   A   B1    Y   VDD   PMOS_3P3   W=Wp  L=0.35um

* X3 Y  Y_inv VDD GND cmos_inv

* CL   Y_inv    GND   cf
VDD  VDD    GND   dd
VGND GND    0     0
.param start=20.0ns delta=0.01ns end=40.0ns
VA0    A0   GND   PWL(0ns 0V `start-delta` 0V start dd `end-delta` dd end 0V)
VB0    B0   GND   PWL(0ns 0V `start-delta` 0V start 0V `end-delta` 0V end 0V)  


.MEASURE TRAN vomax MAX V(Y_inv) FROM 10n TO 20n
.MEASURE TRAN vomin MIN V(Y_inv) FROM 20n TO 30n
.MEASURE TRAN tPHL TRIG V(A) VAL=0.5*dd RISE=1 TARG V(Y) VAL='0.5*(vomax+vomin)' FALL=1
.MEASURE TRAN tPLH TRIG V(B) VAL=0.5*dd FALL=1 TARG V(Y) VAL='0.5*(vomax+vomin)' RISE=2
.MEASURE tran tr TRIG V(Y)='0.1*(vomax-vomin)+vomin' RISE=1 TARG V(Y)='0.9*(vomax-vomin)+vomin' RISE=1
.MEASURE tran tf TRIG V(Y)='0.9*(vomax-vomin)+vomin' FALL=1 TARG V(Y)='0.1*(vomax-vomin)+vomin' FALL=1
.MEASURE tran avgPower AVG P(VDD) FROM=20ns TO=60ns

.tran  0.01ns   100nS 
.probe V(Y) p(VDD) 
**********************************
.END